LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY operative IS
  PORT (

  );
END operative;

ARCHITECTURE operative_arch OF operative IS

  SIGNAL

BEGIN

END ARCHITECTURE operative_arch;
